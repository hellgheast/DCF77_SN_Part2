-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Concurrent Statement 'concurrent0' in architecture 'Behavioral' of entity 'kcpsm3_int_test'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface signals:
-- 
-- in_port : out    std_logic_vector(7 downto 0);
-- reset   : out    std_logic;
-- 
-- EASE/HDL end ----------------------------------------------------------------
in_port <= "00000000";
reset <= '0';
