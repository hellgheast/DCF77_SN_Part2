-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'rtl' of entity 'inversor'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture rtl of inversor is

begin

end architecture rtl ; -- of inversor

