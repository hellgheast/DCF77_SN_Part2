-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'rtl' of entity 'DecodeAdress'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
--   port (
--     adress              : in     std_logic_vector(7 downto 0);
--     adress_dcf          : out    std_logic_vector(3 downto 0);
--     adress_displayblock : out    std_logic_vector(2 downto 0);
--     adress_mux_dcf_test : out    std_logic;
--     dcf_cs              : out    std_logic;
--     displayblock_cs     : out    std_logic;
--     uart_tx_cs          : out    std_logic;
--     write_strobe        : in     std_logic);
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture rtl of DecodeAdress is

begin

end architecture rtl ; -- of DecodeAdress

